ENTITY first_entity IS
    Generic declarations
    Port declarations
END ENTITY;