COMPONENT <lower-level-design-name>
PORT(
    <port_name>:<port_type> <data_type>;
    <port_name>:<port_type> <data_type>;
);
END COMPONENT;