<instance_name> : <lower_level_design_name>
PORT MAP(
    <lower_level_port_name> => <current_level_port_name>,
    <lower_level_port_name> => <current_level_port_name> 
)

[
{question:1, choice:3},
{question:2, choice:2},
{question:3, answer:'Cldl'}
]